LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decoder IS
    PORT ( w  : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
           En : IN  STD_LOGIC;
           y  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) );
END decoder;

ARCHITECTURE Behavior OF decoder IS
    SIGNAL Enw : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
    Enw <= En & w;
    WITH Enw SELECT
        y <= "00000001" WHEN "1000",  -- Enable = 1 and w = 000 (s0)
             "00000010" WHEN "1001",  -- Enable = 1 and w = 001 (s1)
             "00000100" WHEN "1010",  -- Enable = 1 and w = 010 (s2)
             "00001000" WHEN "1011",  -- Enable = 1 and w = 011 (s3)
             "00010000" WHEN "1100",  -- Enable = 1 and w = 100 (s4)
             "00100000" WHEN "1101",  -- Enable = 1 and w = 101 (s5)
             "01000000" WHEN "1110",  -- Enable = 1 and w = 110 (s6)
             "10000000" WHEN "1111",  -- Enable = 1 and w = 111 (s7)
             "00000000" WHEN OTHERS;  -- Default (disabled or invalid inputs)
END Behavior;

